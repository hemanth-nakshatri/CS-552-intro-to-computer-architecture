module ReadDecoder_4_16(Wordline, RegId);
  input [3:0] RegId;
  output [15:0] Wordline;

  assign Wordline = (RegId == 0) ? 16'b0000000000000001 :
                    (RegId == 1) ? 16'b0000000000000010 :
                    (RegId == 2) ? 16'b0000000000000100 :
                    (RegId == 3) ? 16'b0000000000001000 :
                    (RegId == 4) ? 16'b0000000000010000 :
                    (RegId == 5) ? 16'b0000000000100000 :
                    (RegId == 6) ? 16'b0000000001000000 :
                    (RegId == 7) ? 16'b0000000010000000 :
                    (RegId == 8) ? 16'b0000000100000000 :
                    (RegId == 9) ? 16'b0000001000000000 :
                    (RegId == 10) ? 16'b0000010000000000 :
                    (RegId == 11) ? 16'b0000100000000000 :
                    (RegId == 12) ? 16'b0001000000000000 :
                    (RegId == 13) ? 16'b0010000000000000 :
                    (RegId == 14) ? 16'b0100000000000000 :
                    (RegId == 15) ? 16'b1000000000000000 : 16'b0000000000000000;
endmodule

